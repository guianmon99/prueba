----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.05.2022 16:10:42
-- Design Name: 
-- Module Name: 7_seg - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity 7_seg is
    Port ( b : in STD_LOGIC_VECTOR (2 downto 0);
           anode : in STD_LOGIC_VECTOR (3 downto 0);
           catode : in STD_LOGIC_VECTOR (7 downto 0));
end 7_seg;

architecture Behavioral of 7_seg is

begin


end Behavioral;
